entity HelloWorldTb is
end entity;

architecture sim of HelloWorld is begin

    process is begin
        

    end process;

end architecture;